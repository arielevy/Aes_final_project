library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity Inv_Sbox8 is
port(
Data_IN :in std_logic_vector (7 downto 0); -- Data in
Clock : in std_logic; --Clock in
reset : in std_logic;
Data_OUT : out std_logic_vector (7 downto 0) --Data out
);
end Inv_SBox8;

architecture Behav of Inv_SBox8 is

begin
process(Data_IN,clock,reset)	
begin
if (reset = '1') then Data_OUT<=x"00";

elsif (clock'event and clock ='1') then

case Data_IN is -- make look up table
		when x"00" => Data_OUT <= x"52";
		when x"01" => Data_OUT <= x"09";
		when x"02" => Data_OUT <= x"6a";
		when x"03" => Data_OUT <= x"d5";
		when x"04" => Data_OUT <= x"30";
		when x"05" => Data_OUT <= x"36";
		when x"06" => Data_OUT <= x"a5";
		when x"07" => Data_OUT <= x"38";
		when x"08" => Data_OUT <= x"bf";
		when x"09" => Data_OUT <= x"40";
		when x"0a" => Data_OUT <= x"a3";
		when x"0b" => Data_OUT <= x"9e";
		when x"0c" => Data_OUT <= x"81";
		when x"0d" => Data_OUT <= x"f3";
		when x"0e" => Data_OUT <= x"d7";
		when x"0f" => Data_OUT <= x"fb";
		when x"10" => Data_OUT <= x"7c";
		when x"11" => Data_OUT <= x"e3";
		when x"12" => Data_OUT <= x"39";
		when x"13" => Data_OUT <= x"82";
		when x"14" => Data_OUT <= x"9b";
		when x"15" => Data_OUT <= x"2f";
		when x"16" => Data_OUT <= x"ff";
		when x"17" => Data_OUT <= x"87";
		when x"18" => Data_OUT <= x"34";
		when x"19" => Data_OUT <= x"8e";
		when x"1a" => Data_OUT <= x"43";
		when x"1b" => Data_OUT <= x"44";
		when x"1c" => Data_OUT <= x"c4";
		when x"1d" => Data_OUT <= x"de";
		when x"1e" => Data_OUT <= x"e9";
		when x"1f" => Data_OUT <= x"cb";
		when x"20" => Data_OUT <= x"54";
		when x"21" => Data_OUT <= x"7b";
		when x"22" => Data_OUT <= x"94";
		when x"23" => Data_OUT <= x"32";
		when x"24" => Data_OUT <= x"a6";
		when x"25" => Data_OUT <= x"c2";
		when x"26" => Data_OUT <= x"23";
		when x"27" => Data_OUT <= x"3d";
		when x"28" => Data_OUT <= x"ee";
		when x"29" => Data_OUT <= x"4c";
		when x"2a" => Data_OUT <= x"95";
		when x"2b" => Data_OUT <= x"0b";
		when x"2c" => Data_OUT <= x"42";
		when x"2d" => Data_OUT <= x"fa";
		when x"2e" => Data_OUT <= x"c3";
		when x"2f" => Data_OUT <= x"4e";
		when x"30" => Data_OUT <= x"08";
		when x"31" => Data_OUT <= x"2e";
		when x"32" => Data_OUT <= x"a1";
		when x"33" => Data_OUT <= x"66";
		when x"34" => Data_OUT <= x"28";
		when x"35" => Data_OUT <= x"d9";
		when x"36" => Data_OUT <= x"24";
		when x"37" => Data_OUT <= x"b2";
		when x"38" => Data_OUT <= x"76";
		when x"39" => Data_OUT <= x"5b";
		when x"3a" => Data_OUT <= x"a2";
		when x"3b" => Data_OUT <= x"49";
		when x"3c" => Data_OUT <= x"6d";
		when x"3d" => Data_OUT <= x"8b";
		when x"3e" => Data_OUT <= x"d1";
		when x"3f" => Data_OUT <= x"25";
		when x"40" => Data_OUT <= x"72";
		when x"41" => Data_OUT <= x"f8";
		when x"42" => Data_OUT <= x"f6";
		when x"43" => Data_OUT <= x"64";
		when x"44" => Data_OUT <= x"86";
		when x"45" => Data_OUT <= x"68";
		when x"46" => Data_OUT <= x"98";
		when x"47" => Data_OUT <= x"16";
		when x"48" => Data_OUT <= x"d4";
		when x"49" => Data_OUT <= x"a4";
		when x"4a" => Data_OUT <= x"5c";
		when x"4b" => Data_OUT <= x"cc";
		when x"4c" => Data_OUT <= x"5d";
		when x"4d" => Data_OUT <= x"65";
		when x"4e" => Data_OUT <= x"b6";
		when x"4f" => Data_OUT <= x"92";
		when x"50" => Data_OUT <= x"6c";
		when x"51" => Data_OUT <= x"70";
		when x"52" => Data_OUT <= x"48";
		when x"53" => Data_OUT <= x"50";
		when x"54" => Data_OUT <= x"fd";
		when x"55" => Data_OUT <= x"ed";
		when x"56" => Data_OUT <= x"b9";
		when x"57" => Data_OUT <= x"da";
		when x"58" => Data_OUT <= x"5e";
		when x"59" => Data_OUT <= x"15";
		when x"5a" => Data_OUT <= x"46";
		when x"5b" => Data_OUT <= x"57";
		when x"5c" => Data_OUT <= x"a7";
		when x"5d" => Data_OUT <= x"8d";
		when x"5e" => Data_OUT <= x"9d";
		when x"5f" => Data_OUT <= x"84";
		when x"60" => Data_OUT <= x"90";
		when x"61" => Data_OUT <= x"d8";
		when x"62" => Data_OUT <= x"ab";
		when x"63" => Data_OUT <= x"00";
		when x"64" => Data_OUT <= x"8c";
		when x"65" => Data_OUT <= x"bc";
		when x"66" => Data_OUT <= x"d3";
		when x"67" => Data_OUT <= x"0a";
		when x"68" => Data_OUT <= x"f7";
		when x"69" => Data_OUT <= x"e4";
		when x"6a" => Data_OUT <= x"58";
		when x"6b" => Data_OUT <= x"05";
		when x"6c" => Data_OUT <= x"b8";
		when x"6d" => Data_OUT <= x"b3";
		when x"6e" => Data_OUT <= x"45";
		when x"6f" => Data_OUT <= x"06";
		when x"70" => Data_OUT <= x"d0";
		when x"71" => Data_OUT <= x"2c";
		when x"72" => Data_OUT <= x"1e";
		when x"73" => Data_OUT <= x"8f";
		when x"74" => Data_OUT <= x"ca";
		when x"75" => Data_OUT <= x"3f";
		when x"76" => Data_OUT <= x"0f";
		when x"77" => Data_OUT <= x"02";
		when x"78" => Data_OUT <= x"c1";
		when x"79" => Data_OUT <= x"af";
		when x"7a" => Data_OUT <= x"bd";
		when x"7b" => Data_OUT <= x"03";
		when x"7c" => Data_OUT <= x"01";
		when x"7d" => Data_OUT <= x"13";
		when x"7e" => Data_OUT <= x"8a";
		when x"7f" => Data_OUT <= x"6b";
		when x"80" => Data_OUT <= x"3a";
		when x"81" => Data_OUT <= x"91";
		when x"82" => Data_OUT <= x"11";
		when x"83" => Data_OUT <= x"41";
		when x"84" => Data_OUT <= x"4f";
		when x"85" => Data_OUT <= x"67";
		when x"86" => Data_OUT <= x"dc";
		when x"87" => Data_OUT <= x"ea";
		when x"88" => Data_OUT <= x"97";
		when x"89" => Data_OUT <= x"f2";
		when x"8a" => Data_OUT <= x"cf";
		when x"8b" => Data_OUT <= x"ce";
		when x"8c" => Data_OUT <= x"f0";
		when x"8d" => Data_OUT <= x"b4";
		when x"8e" => Data_OUT <= x"e6";
		when x"8f" => Data_OUT <= x"73";
		when x"90" => Data_OUT <= x"96";
		when x"91" => Data_OUT <= x"ac";
		when x"92" => Data_OUT <= x"74";
		when x"93" => Data_OUT <= x"22";
		when x"94" => Data_OUT <= x"e7";
		when x"95" => Data_OUT <= x"ad";
		when x"96" => Data_OUT <= x"35";
		when x"97" => Data_OUT <= x"85";
		when x"98" => Data_OUT <= x"e2";
		when x"99" => Data_OUT <= x"f9";
		when x"9a" => Data_OUT <= x"37";
		when x"9b" => Data_OUT <= x"e8";
		when x"9c" => Data_OUT <= x"1c";
		when x"9d" => Data_OUT <= x"75";
		when x"9e" => Data_OUT <= x"df";
		when x"9f" => Data_OUT <= x"6e";
		when x"a0" => Data_OUT <= x"47";
		when x"a1" => Data_OUT <= x"f1";
		when x"a2" => Data_OUT <= x"1a";
		when x"a3" => Data_OUT <= x"71";
		when x"a4" => Data_OUT <= x"1d";
		when x"a5" => Data_OUT <= x"29";
		when x"a6" => Data_OUT <= x"c5";
		when x"a7" => Data_OUT <= x"89";
		when x"a8" => Data_OUT <= x"6f";
		when x"a9" => Data_OUT <= x"b7";
		when x"aa" => Data_OUT <= x"62";
		when x"ab" => Data_OUT <= x"0e";
		when x"ac" => Data_OUT <= x"aa";
		when x"ad" => Data_OUT <= x"18";
		when x"ae" => Data_OUT <= x"be";
		when x"af" => Data_OUT <= x"1b";
		when x"b0" => Data_OUT <= x"fc";
		when x"b1" => Data_OUT <= x"56";
		when x"b2" => Data_OUT <= x"3e";
		when x"b3" => Data_OUT <= x"4b";
		when x"b4" => Data_OUT <= x"c6";
		when x"b5" => Data_OUT <= x"d2";
		when x"b6" => Data_OUT <= x"79";
		when x"b7" => Data_OUT <= x"20";
		when x"b8" => Data_OUT <= x"9a";
		when x"b9" => Data_OUT <= x"db";
		when x"ba" => Data_OUT <= x"c0";
		when x"bb" => Data_OUT <= x"fe";
		when x"bc" => Data_OUT <= x"78";
		when x"bd" => Data_OUT <= x"cd";
		when x"be" => Data_OUT <= x"5a";
		when x"bf" => Data_OUT <= x"f4";
		when x"c0" => Data_OUT <= x"1f";
		when x"c1" => Data_OUT <= x"dd";
		when x"c2" => Data_OUT <= x"a8";
		when x"c3" => Data_OUT <= x"33";
		when x"c4" => Data_OUT <= x"88";
		when x"c5" => Data_OUT <= x"07";
		when x"c6" => Data_OUT <= x"c7";
		when x"c7" => Data_OUT <= x"31";
		when x"c8" => Data_OUT <= x"b1";
		when x"c9" => Data_OUT <= x"12";
		when x"ca" => Data_OUT <= x"10";
		when x"cb" => Data_OUT <= x"59";
		when x"cc" => Data_OUT <= x"27";
		when x"cd" => Data_OUT <= x"80";
		when x"ce" => Data_OUT <= x"ec";
		when x"cf" => Data_OUT <= x"5f";
		when x"d0" => Data_OUT <= x"60";
		when x"d1" => Data_OUT <= x"51";
		when x"d2" => Data_OUT <= x"7f";
		when x"d3" => Data_OUT <= x"a9";
		when x"d4" => Data_OUT <= x"19";
		when x"d5" => Data_OUT <= x"b5";
		when x"d6" => Data_OUT <= x"4a";
		when x"d7" => Data_OUT <= x"0d";
		when x"d8" => Data_OUT <= x"2d";
		when x"d9" => Data_OUT <= x"e5";
		when x"da" => Data_OUT <= x"7a";
		when x"db" => Data_OUT <= x"9f";
		when x"dc" => Data_OUT <= x"93";
		when x"dd" => Data_OUT <= x"c9";
		when x"de" => Data_OUT <= x"9c";
		when x"df" => Data_OUT <= x"ef";
		when x"e0" => Data_OUT <= x"a0";
		when x"e1" => Data_OUT <= x"e0";
		when x"e2" => Data_OUT <= x"3b";
		when x"e3" => Data_OUT <= x"4d";
		when x"e4" => Data_OUT <= x"ae";
		when x"e5" => Data_OUT <= x"2a";
		when x"e6" => Data_OUT <= x"f5";
		when x"e7" => Data_OUT <= x"b0";
		when x"e8" => Data_OUT <= x"c8";
		when x"e9" => Data_OUT <= x"eb";
		when x"ea" => Data_OUT <= x"bb";
		when x"eb" => Data_OUT <= x"3c";
		when x"ec" => Data_OUT <= x"83";
		when x"ed" => Data_OUT <= x"53";
		when x"ee" => Data_OUT <= x"99";
		when x"ef" => Data_OUT <= x"61";
		when x"f0" => Data_OUT <= x"17";
		when x"f1" => Data_OUT <= x"2b";
		when x"f2" => Data_OUT <= x"04";
		when x"f3" => Data_OUT <= x"7e";
		when x"f4" => Data_OUT <= x"ba";
		when x"f5" => Data_OUT <= x"77";
		when x"f6" => Data_OUT <= x"d6";
		when x"f7" => Data_OUT <= x"26";
		when x"f8" => Data_OUT <= x"e1";
		when x"f9" => Data_OUT <= x"69";
		when x"fa" => Data_OUT <= x"14";
		when x"fb" => Data_OUT <= x"63";
		when x"fc" => Data_OUT <= x"55";
		when x"fd" => Data_OUT <= x"21";
		when x"fe" => Data_OUT <= x"0c";
		when x"ff" => Data_OUT <= x"7d";
			when others=> Data_OUT<=x"52";
end case;

end if;		
end process;
end architecture;