library ieee;
use ieee.std_logic_1164.all;
use ieee.std_logic_unsigned.all;

entity Sbox8 is
port(
Data_IN :in std_logic_vector (7 downto 0); -- Data in
Clock : in std_logic; --Clock in
reset : in std_logic;
Data_OUT : out std_logic_vector (7 downto 0) --Data out
);
end SBox8;

architecture Behav of SBox8 is

begin
process(Data_IN,clock,reset)	
begin
if (reset = '1') then Data_OUT<=x"00";

elsif (clock'event and clock ='1') then

case Data_IN is -- make lookup table
			when "00000000"=>Data_OUT<=x"63";
			when "00000001"=>Data_OUT<=x"7c";
			when "00000010"=>Data_OUT<=x"77";
			when "00000011"=>Data_OUT<=x"7b";
			when "00000100"=>Data_OUT<=x"f2";
			when "00000101"=>Data_OUT<=x"6b";
			when "00000110"=>Data_OUT<=x"6f";
			when "00000111"=>Data_OUT<=x"c5";
			when "00001000"=>Data_OUT<=x"30";
			when "00001001"=>Data_OUT<=x"01";
			when "00001010"=>Data_OUT<=x"67";
			when "00001011"=>Data_OUT<=x"2b";
			when "00001100"=>Data_OUT<=x"fe";
			when "00001101"=>Data_OUT<=x"d7";
			when "00001110"=>Data_OUT<=x"ab";
			when "00001111"=>Data_OUT<=x"76";
			when "00010000"=>Data_OUT<=x"ca";
			when "00010001"=>Data_OUT<=x"82";
			when "00010010"=>Data_OUT<=x"c9";
			when "00010011"=>Data_OUT<=x"7d";
			when "00010100"=>Data_OUT<=x"fa";
			when "00010101"=>Data_OUT<=x"59";
			when "00010110"=>Data_OUT<=x"47";
			when "00010111"=>Data_OUT<=x"f0";
			when "00011000"=>Data_OUT<=x"ad";
			when "00011001"=>Data_OUT<=x"d4";
			when "00011010"=>Data_OUT<=x"a2";
			when "00011011"=>Data_OUT<=x"af";
			when "00011100"=>Data_OUT<=x"9c";
			when "00011101"=>Data_OUT<=x"a4";
			when "00011110"=>Data_OUT<=x"72";
			when "00011111"=>Data_OUT<=x"c0";
			when "00100000"=>Data_OUT<=x"b7";
			when "00100001"=>Data_OUT<=x"fd";
			when "00100010"=>Data_OUT<=x"93";
			when "00100011"=>Data_OUT<=x"26";
			when "00100100"=>Data_OUT<=x"36";
			when "00100101"=>Data_OUT<=x"3f";
			when "00100110"=>Data_OUT<=x"f7";
			when "00100111"=>Data_OUT<=x"cc";
			when "00101000"=>Data_OUT<=x"34";
			when "00101001"=>Data_OUT<=x"a5";
			when "00101010"=>Data_OUT<=x"e5";
			when "00101011"=>Data_OUT<=x"f1";
			when "00101100"=>Data_OUT<=x"71";
			when "00101101"=>Data_OUT<=x"d8";
			when "00101110"=>Data_OUT<=x"31";
			when "00101111"=>Data_OUT<=x"15";
			when "00110000"=>Data_OUT<=x"04";
			when "00110001"=>Data_OUT<=x"c7";
			when "00110010"=>Data_OUT<=x"23";
			when "00110011"=>Data_OUT<=x"c3";
			when "00110100"=>Data_OUT<=x"18";
			when "00110101"=>Data_OUT<=x"96";				
			when "00110110"=>Data_OUT<=x"05";
			when "00110111"=>Data_OUT<=x"9a";
			when "00111000"=>Data_OUT<=x"07";
			when "00111001"=>Data_OUT<=x"12";
			when "00111010"=>Data_OUT<=x"80";
			when "00111011"=>Data_OUT<=x"e2";
			when "00111100"=>Data_OUT<=x"eb";
			when "00111101"=>Data_OUT<=x"27";
			when "00111110"=>Data_OUT<=x"b2";
			when "00111111"=>Data_OUT<=x"75";
			when "01000000"=>Data_OUT<=x"09";
			when "01000001"=>Data_OUT<=x"83";
			when "01000010"=>Data_OUT<=x"2c";
			when "01000011"=>Data_OUT<=x"1a";
			when "01000100"=>Data_OUT<=x"1b";
			when "01000101"=>Data_OUT<=x"6e";
			when "01000110"=>Data_OUT<=x"5a";
         when "01000111"=>Data_OUT<=x"a0";
			when "01001000"=>Data_OUT<=x"52";
			when "01001001"=>Data_OUT<=x"3b";
			when "01001010"=>Data_OUT<=x"d6";
			when "01001011"=>Data_OUT<=x"b3";
			when "01001100"=>Data_OUT<=x"29";
			when "01001101"=>Data_OUT<=x"e3";
			when "01001110"=>Data_OUT<=x"2f";
		   when "01001111"=>Data_OUT<=x"84";
			when "01010000"=>Data_OUT<=x"53";
			when "01010001"=>Data_OUT<=x"d1";
			when "01010010"=>Data_OUT<=x"00";
			when "01010011"=>Data_OUT<=x"ed";
			when "01010100"=>Data_OUT<=x"20";
			when "01010101"=>Data_OUT<=x"fc";
			when "01010110"=>Data_OUT<=x"b1";
			when "01010111"=>Data_OUT<=x"5b";
			when "01011000"=>Data_OUT<=x"6a";
			when "01011001"=>Data_OUT<=x"cb";
			when "01011010"=>Data_OUT<=x"be";
			when "01011011"=>Data_OUT<=x"39";
			when "01011100"=>Data_OUT<=x"4a";
			when "01011101"=>Data_OUT<=x"4c";
			when "01011110"=>Data_OUT<=x"58";
			when "01011111"=>Data_OUT<=x"cf";
			when "01100000"=>Data_OUT<=x"d0";
			when "01100001"=>Data_OUT<=x"ef";
			when "01100010"=>Data_OUT<=x"aa";
			when "01100011"=>Data_OUT<=x"fb";
			when "01100100"=>Data_OUT<=x"43";
			when "01100101"=>Data_OUT<=x"4d";
			when "01100110"=>Data_OUT<=x"33";
			when "01100111"=>Data_OUT<=x"85";
			when "01101000"=>Data_OUT<=x"45";
			when "01101001"=>Data_OUT<=x"f9";
		   when "01101010"=>Data_OUT<=x"02";
			when "01101011"=>Data_OUT<=x"7f";
			when "01101100"=>Data_OUT<=x"50";
			when "01101101"=>Data_OUT<=x"3c";
			when "01101110"=>Data_OUT<=x"9f";
			when "01101111"=>Data_OUT<=x"a8";
			when "01110000"=>Data_OUT<=x"51";
			when "01110001"=>Data_OUT<=x"a3";
			when "01110010"=>Data_OUT<=x"40";
			when "01110011"=>Data_OUT<=x"8f";
			when "01110100"=>Data_OUT<=x"92";
			when "01110101"=>Data_OUT<=x"9d";
			when "01110110"=>Data_OUT<=x"38";
		   when "01110111"=>Data_OUT<=x"f5";
			when "01111000"=>Data_OUT<=x"bc";
			when "01111001"=>Data_OUT<=x"b6";
			when "01111010"=>Data_OUT<=x"da";
			when "01111011"=>Data_OUT<=x"21";
			when "01111100"=>Data_OUT<=x"10";
			when "01111101"=>Data_OUT<=x"ff";
			when "01111110"=>Data_OUT<=x"f3";
			when "01111111"=>Data_OUT<=x"d2";
			when "10000000"=>Data_OUT<=x"cd";
			when "10000001"=>Data_OUT<=x"0c";
			when "10000010"=>Data_OUT<=x"13";
			when "10000011"=>Data_OUT<=x"ec";
			when "10000100"=>Data_OUT<=x"5f";
			when "10000101"=>Data_OUT<=x"97";
			when "10000110"=>Data_OUT<=x"44";
			when "10000111"=>Data_OUT<=x"17";
			when "10001000"=>Data_OUT<=x"c4";
			when "10001001"=>Data_OUT<=x"a7";
			when "10001010"=>Data_OUT<=x"7e";
			when "10001011"=>Data_OUT<=x"3d";
			when "10001100"=>Data_OUT<=x"64";
			when "10001101"=>Data_OUT<=x"5d";
			when "10001110"=>Data_OUT<=x"19";
			when "10001111"=>Data_OUT<=x"73";
			when "10010000"=>Data_OUT<=x"60";
			when "10010001"=>Data_OUT<=x"81";
			when "10010010"=>Data_OUT<=x"4f";
			when "10010011"=>Data_OUT<=x"dc";
			when "10010100"=>Data_OUT<=x"22";
			when "10010101"=>Data_OUT<=x"2a";
			when "10010110"=>Data_OUT<=x"90";
			when "10010111"=>Data_OUT<=x"88";
			when "10011000"=>Data_OUT<=x"46";
			when "10011001"=>Data_OUT<=x"ee";
			when "10011010"=>Data_OUT<=x"b8";
			when "10011011"=>Data_OUT<=x"14";
			when "10011100"=>Data_OUT<=x"de";
			when "10011101"=>Data_OUT<=x"5e";
			when "10011110"=>Data_OUT<=x"0b";
			when "10011111"=>Data_OUT<=x"db";
			when "10100000"=>Data_OUT<=x"e0";
			when "10100001"=>Data_OUT<=x"32";
			when "10100010"=>Data_OUT<=x"3a";
			when "10100011"=>Data_OUT<=x"0a";
			when "10100100"=>Data_OUT<=x"49";
			when "10100101"=>Data_OUT<=x"06";
			when "10100110"=>Data_OUT<=x"24";
			when "10100111"=>Data_OUT<=x"5c";
			when "10101000"=>Data_OUT<=x"c2";
			when "10101001"=>Data_OUT<=x"d3";
			when "10101010"=>Data_OUT<=x"ac";
			when "10101011"=>Data_OUT<=x"62";
			when "10101100"=>Data_OUT<=x"91";
			when "10101101"=>Data_OUT<=x"95";
			when "10101110"=>Data_OUT<=x"e4";
			when "10101111"=>Data_OUT<=x"79";
			when "10110000"=>Data_OUT<=x"e7";
			when "10110001"=>Data_OUT<=x"c8";
			when "10110010"=>Data_OUT<=x"37";
			when "10110011"=>Data_OUT<=x"6d";
			when "10110100"=>Data_OUT<=x"8d";
			when "10110101"=>Data_OUT<=x"d5";
			when "10110110"=>Data_OUT<=x"4e";
			when "10110111"=>Data_OUT<=x"a9";
			when "10111000"=>Data_OUT<=x"6c";
			when "10111001"=>Data_OUT<=x"56";
			when "10111010"=>Data_OUT<=x"f4";
			when "10111011"=>Data_OUT<=x"ea";
			when "10111100"=>Data_OUT<=x"65";
			when "10111101"=>Data_OUT<=x"7a";
			when "10111110"=>Data_OUT<=x"ae";
			when "10111111"=>Data_OUT<=x"08";
			when "11000000"=>Data_OUT<=x"ba";
			when "11000001"=>Data_OUT<=x"78";
			when "11000010"=>Data_OUT<=x"25";
			when "11000011"=>Data_OUT<=x"2e";
			when "11000100"=>Data_OUT<=x"1c";
			when "11000101"=>Data_OUT<=x"a6";
			when "11000110"=>Data_OUT<=x"b4";
			when "11000111"=>Data_OUT<=x"c6";
			when "11001000"=>Data_OUT<=x"e8";
			when "11001001"=>Data_OUT<=x"dd";
			when "11001010"=>Data_OUT<=x"74";
			when "11001011"=>Data_OUT<=x"1f";
			when "11001100"=>Data_OUT<=x"4b";
			when "11001101"=>Data_OUT<=x"bd";
			when "11001110"=>Data_OUT<=x"8b";
			when "11001111"=>Data_OUT<=x"8a";
			when "11010000"=>Data_OUT<=x"70";
			when "11010001"=>Data_OUT<=x"3e";
			when "11010010"=>Data_OUT<=x"b5";
			when "11010011"=>Data_OUT<=x"66";
			when "11010100"=>Data_OUT<=x"48";
			when "11010101"=>Data_OUT<=x"03";
			when "11010110"=>Data_OUT<=x"f6";
		   when "11010111"=>Data_OUT<=x"0e";
			when "11011000"=>Data_OUT<=x"61";
			when "11011001"=>Data_OUT<=x"35";
			when "11011010"=>Data_OUT<=x"57";
			when "11011011"=>Data_OUT<=x"b9";
			when "11011100"=>Data_OUT<=x"86";
			when "11011101"=>Data_OUT<=x"c1";
			when "11011110"=>Data_OUT<=x"1d";
			when "11011111"=>Data_OUT<=x"9e";
			when "11100000"=>Data_OUT<=x"e1";
			when "11100001"=>Data_OUT<=x"f8";
			when "11100010"=>Data_OUT<=x"98";
			when "11100011"=>Data_OUT<=x"11";
			when "11100100"=>Data_OUT<=x"69";
			when "11100101"=>Data_OUT<=x"d9";
			when "11100110"=>Data_OUT<=x"8e";
			when "11100111"=>Data_OUT<=x"94";
			when "11101000"=>Data_OUT<=x"9b";
			when "11101001"=>Data_OUT<=x"1e";
			when "11101010"=>Data_OUT<=x"87";
			when "11101011"=>Data_OUT<=x"e9";
			when "11101100"=>Data_OUT<=x"ce";
			when "11101101"=>Data_OUT<=x"55";
			when "11101110"=>Data_OUT<=x"28";
			when "11101111"=>Data_OUT<=x"df";
			when "11110000"=>Data_OUT<=x"8c";
			when "11110001"=>Data_OUT<=x"a1";
			when "11110010"=>Data_OUT<=x"89";
			when "11110011"=>Data_OUT<=x"0d";
			when "11110100"=>Data_OUT<=x"bf";
			when "11110101"=>Data_OUT<=x"e6";
			when "11110110"=>Data_OUT<=x"42";
			when "11110111"=>Data_OUT<=x"68";
			when "11111000"=>Data_OUT<=x"41";
			when "11111001"=>Data_OUT<=x"99";
			when "11111010"=>Data_OUT<=x"2d";
			when "11111011"=>Data_OUT<=x"0f";
			when "11111100"=>Data_OUT<=x"b0";
			when "11111101"=>Data_OUT<=x"54";
			when "11111110"=>Data_OUT<=x"bb";
			when others=> Data_OUT<=x"16";
end case;

end if;		
end process;
end architecture;